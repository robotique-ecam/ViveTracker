`define F_1MHz 12
`define F_2MHz 6
`define F_3MHz 4
`define F_4MHz 3

`define F_1KHz 12_000
`define F_2KHz 6_000
`define F_3KHz 4_000
`define F_4KHz 3_000

`define F_4Hz 3_000_000
`define F_3Hz 4_000_000
`define F_2Hz 6_000_000
`define F_1Hz 12_000_000
